module IFetcher(
input logic clk,
input logic[31:0] PC,
output logic[63:0] instruction_o
);


endmodule