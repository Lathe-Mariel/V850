module Writeback(

);


endmodule