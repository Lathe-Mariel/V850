module Memory(

);


endmodule