module adder(
wire clk,
logic[31:0] reg1,
logic[31:0] reg2
);

always @(posedge clk)begin
//    reg1 <= reg1 + reg2;
end

endmodule